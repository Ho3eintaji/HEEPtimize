// Copyright 2022 EPFL and Politecnico di Torino.
// Solderpad Hardware License, Version 2.1, see LICENSE.md for details.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// File: pad_cell_input.sv
// Author: Michele Caon
// Date: 14/05/2023
// Description: Inpud pad standard cell

module pad_cell_input #(
  parameter int unsigned PADATTR = 16
) (
  input logic pad_in_i, // pad input value
  input logic pad_oe_i, // pad output enable
  output logic pad_out_o, // pad output value
  input logic pad_io, // pad value
  input logic [PADATTR-1:0] pad_attributes_i // pad attributes
);
  // TSMC65 pad standard cell
  tsmc65_pad_cell_input #(
    .PADATTR (PADATTR )
  ) u_pad_cell_input (
  	.pad_in_i         (pad_in_i         ),
    .pad_oe_i         (pad_oe_i         ),
    .pad_out_o        (pad_out_o        ),
    .pad_io           (pad_io           ),
    .pad_attributes_i (pad_attributes_i )
  );
endmodule
